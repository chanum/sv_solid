
class base_transaction;
  // common properties and methods
endclass

class extended_transaction extends base_transaction;
  // additional properties and methods
endclass