
module counter #(parameter WIDTH = 8) (
  input logic   clk,
  input logic   reset,
  output logic  [WIDTH-1:0] count_o
);

  // counter implementation

endmodule : counter
