class base_transaction;
  // Propiedades y métodos comunes
endclass

class extended_transaction extends base_transaction;
  // Propiedades y métodos adicionales
endclass